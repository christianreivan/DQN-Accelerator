module Action_determiner (
    clk, rst, step, controller, episode,
    Qst_0, Qst_1, Qst_2, Qst_3, 
    Qst1_0, Qst1_1, Qst1_2, Qst1_3, act, st, st1, Qt, maxQt1
);

    input clk, rst;
    input [3:0] step, controller;
    input [11:0] episode;
    input [15:0] Qst_0, Qst_1, Qst_2, Qst_3;
    input [15:0] Qst1_0, Qst1_1, Qst1_2, Qst1_3;
    output [1:0] act;
    output [3:0] st, st1;
    output [15:0] Qt, maxQt1;

    wire comparison_result;
    wire [1:0] qmax_act, random_act;

    qnext_max qnex_max_mod(
        Qst1_0, Qst1_1, Qst1_2, Qst1_3, maxQt1
    );
    qmax_action qmaxact_mod(
        Qst_0, Qst_1, Qst_2, Qst_3, Qt, qmax_act
    );
    random_action randomact_mod(
        clk, episode, random_act, comparison_result
    );

    assign act = comparison_result? qmax_act : random_act;

    checker check(
        clk, rst, act, step, controller, st, st1
    );

endmodule
////////////////////////////////////////////////////
//qnext_max
module qnext_max (
    Qst1_0, Qst1_1, Qst1_2, Qst1_3, maxQt1
);
    input signed [15:0] Qst1_0, Qst1_1, Qst1_2, Qst1_3;
    output signed [15:0] maxQt1;

    wire signed [15:0] wire1, wire2;

    assign wire1 = (Qst1_0 > Qst1_1)? Qst1_0 : Qst1_1;
    assign wire2 = (Qst1_2 > Qst1_3)? Qst1_2 : Qst1_3;
    assign maxQt1 = (wire1 > wire2)? wire1 : wire2;
endmodule

////////////////////////////////////////////////////

//qmax_action is a module that generates qmax_action from 
//qvalue generated by neural network
module qmax_action (
    Qst_0, Qst_1, Qst_2, Qst_3, Qt, qmax_act
);
    input signed [15:0] Qst_0, Qst_1, Qst_2, Qst_3;
    output [1:0] qmax_act;
    output signed [15:0] Qt;

    parameter right = 2'd0; 
    parameter up = 2'd1; 
    parameter left = 2'd2; 
    parameter down = 2'd3;

    wire signed [15:0] wire1, wire2, wire3;

    //search the max qvalue
    assign wire1 = (Qst_0 > Qst_1)? Qst_0 : Qst_1;
    assign wire2 = (Qst_2 > Qst_3)? Qst_2 : Qst_3;
    assign wire3 = (wire1 > wire2)? wire1 : wire2;
    
    assign Qt = wire3;
    //qmax action is determined by which qvalue that equal with max qvalue
    assign qmax_act = (wire3 == Qst_0)? right :
                        (wire3 == Qst_1)? up :
                        (wire3 == Qst_2)? left : down;
endmodule

////////////////////////////////////////////////////

//LFSR is a module that generates 12bit random number
module LFSR(clk, random);
    input clk; 
    output [11:0] random; 
    
    reg [11:0] reg_rand; 
    wire feedback; 

    parameter init = 12'b001010010110; 
    initial reg_rand = init; 
    assign feedback = reg_rand[10] ^ reg_rand[7]; 
    
    always @ (posedge clk) begin 
        reg_rand = {reg_rand[10:0], feedback}; 
    end
    
    assign random = reg_rand; 
endmodule

//random_act is a module that generates random_act and comparison of episode-random number
module random_action(
    clk, episode, random_act, comparison_result
);
    input clk;
    input [11:0] episode;
    output comparison_result;
    output [1:0] random_act;

    wire [11:0] random;

    LFSR random_generator(clk, random);

    //if episode < random, the action will be taken is random_act
    //else, the action will be taken is qmax_act
    assign comparison_result = (episode < random)? 1'b1 : 1'b0;

    //assign random_act by taking 2 LSB of random number
    assign random_act = random[1:0];
endmodule

////////////////////////////////////////////////////
module checker (
    clk, rst, act, step, controller, st, st1
);
    input clk, rst;
    input [1:0] act;
    input [3:0] step, controller;
    output [3:0] st, st1;

    reg [3:0] st_temp, st1_temp;
	 
	 assign st = st_temp;
	 assign st1 = st1_temp;
	 
    always @(posedge clk ) begin
        if (rst) 
        begin
            st_temp <= 4'd1;
            st1_temp <= 4'd1;
        end 
        else 
        begin
            if(step != 4'd0) begin
                if(controller == 4'd1)
                 begin
                    st_temp <= st1_temp;
                 end
                else 
                begin
                    if(controller == 4'd6) 
                    begin
                        if (step == 4'd14) begin
                            st1_temp <= 4'd1;
                        end 
                        else 
                        begin
                            
                        end
                        case (act)
                            2'd0 : begin //right
                                if((st_temp == 4'd3) || (st_temp == 4'd6) || (st_temp == 4'd9)) begin
                                    st1_temp <= st_temp;
                                end
                                else  st1_temp <= st_temp + 4'd1;
                            end
                            2'd1 : begin //up
                                if((st_temp == 4'd1) || (st_temp == 4'd2) || (st_temp == 4'd3)) begin
                                    st1_temp <= st_temp;
                                end
                                else  st1_temp <= st_temp - 4'd3;
                            end
                            2'd2 : begin //left
                                if((st_temp == 4'd1) || (st_temp == 4'd4) || (st_temp == 4'd7)) begin
                                    st1_temp <= st_temp;
                                end
                                else  st1_temp <= st_temp - 4'd1;
                            end
                            2'd3 : begin //down
                                if((st_temp == 4'd7) || (st_temp == 4'd8) || (st_temp == 4'd9)) begin
                                    st1_temp <= st_temp;
                                end
                                else  st1_temp <= st_temp + 4'd3;
                            end
                        endcase
                    end
                    else begin
                        st1_temp <= st1_temp;
                        st_temp  <= st_temp;
                    end
                end
            end
            else begin
                st_temp <= st_temp;
                st1_temp <= st1_temp;
            end
        end
    end
endmodule

///////////////////////////////////////////////
///////////////////////////////////////////////

module checker_tb ();
    reg clk, rst;
    reg [1:0] act;
    reg [3:0] step, controller;
    wire [3:0] st, st1;

    checker check_mod(
        clk, rst, act, step, controller, st, st1
    );

    initial begin 
        clk = 1'b1;
        forever #50 clk = ~clk;
    end
    initial begin
        rst = 1;
        act = 2'd0;
    end

endmodule




module regpos (
    clk, rst, controller, din, dout
);
    input clk, rst;
    input [3:0] controller, din;
    output reg [1:0] dout;

    always @(posedge clk ) begin
        if (rst) begin
            dout <= 2'd1;
        end else begin
            if(controller == 4'd1) begin
                dout <= din;    
            end
            else 
                dout <= dout;
        end
    end
endmodule

module regstate (
    clk, rst, controller, din, dout
);
    input clk, rst;
    input [3:0] controller, din;
    output reg [3:0] dout;

    always @(posedge clk ) begin
        if (rst) begin
            dout <= 4'd1;
        end else begin
            if(controller == 4'd1) begin
                dout <= din;    
            end
            else 
                dout <= dout;
        end
    end
endmodule